VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO rom_tvbgone_32k
  CLASS BLOCK ;
  FOREIGN rom_tvbgone_32k ;
  ORIGIN 0.000 0.000 ;
  SIZE 144.900 BY 112.300 ;
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.675000 ;
    PORT
      LAYER met2 ;
        RECT 144.600 8.310 144.900 8.570 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.675000 ;
    PORT
      LAYER met2 ;
        RECT 144.600 9.310 144.900 9.570 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.675000 ;
    PORT
      LAYER met2 ;
        RECT 144.600 10.310 144.900 10.570 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.675000 ;
    PORT
      LAYER met2 ;
        RECT 144.600 11.310 144.900 11.570 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.675000 ;
    PORT
      LAYER met2 ;
        RECT 144.600 12.310 144.900 12.570 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.675000 ;
    PORT
      LAYER met2 ;
        RECT 144.600 7.310 144.900 7.570 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.675000 ;
    PORT
      LAYER met2 ;
        RECT 144.600 6.310 144.900 6.570 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.675000 ;
    PORT
      LAYER met2 ;
        RECT 144.600 5.310 144.900 5.570 ;
    END
  END addr[7]
  PIN addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.675000 ;
    PORT
      LAYER met2 ;
        RECT 144.600 4.310 144.900 4.570 ;
    END
  END addr[8]
  PIN addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.675000 ;
    PORT
      LAYER met2 ;
        RECT 144.600 3.310 144.900 3.570 ;
    END
  END addr[9]
  PIN addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.675000 ;
    PORT
      LAYER met2 ;
        RECT 144.600 2.310 144.900 2.570 ;
    END
  END addr[10]
  PIN addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.675000 ;
    PORT
      LAYER met2 ;
        RECT 144.600 1.310 144.900 1.570 ;
    END
  END addr[11]
  PIN q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.490000 ;
    PORT
      LAYER met2 ;
        RECT 144.600 23.335 144.900 23.595 ;
    END
  END q[0]
  PIN q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.490000 ;
    PORT
      LAYER met2 ;
        RECT 144.600 35.435 144.900 35.695 ;
    END
  END q[1]
  PIN q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.490000 ;
    PORT
      LAYER met2 ;
        RECT 144.600 48.235 144.900 48.495 ;
    END
  END q[2]
  PIN q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.490000 ;
    PORT
      LAYER met2 ;
        RECT 144.600 60.335 144.900 60.595 ;
    END
  END q[3]
  PIN q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.490000 ;
    PORT
      LAYER met2 ;
        RECT 144.600 73.135 144.900 73.395 ;
    END
  END q[4]
  PIN q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.490000 ;
    PORT
      LAYER met2 ;
        RECT 144.600 85.235 144.900 85.495 ;
    END
  END q[5]
  PIN q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.490000 ;
    PORT
      LAYER met2 ;
        RECT 144.600 98.035 144.900 98.295 ;
    END
  END q[6]
  PIN q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.490000 ;
    PORT
      LAYER met2 ;
        RECT 144.600 110.135 144.900 110.395 ;
    END
  END q[7]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.555 10.865 130.285 11.365 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.055 7.445 138.755 8.695 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.755 9.195 137.350 10.445 ;
    END
  END VPWR
  OBS
      LAYER nwell ;
        RECT 0.400 0.000 144.385 112.100 ;
      LAYER li1 ;
        RECT 0.585 0.130 144.295 111.980 ;
      LAYER met1 ;
        RECT 0.055 0.130 144.355 112.115 ;
      LAYER met2 ;
        RECT 0.055 110.675 144.600 111.375 ;
        RECT 0.055 109.855 144.320 110.675 ;
        RECT 0.055 98.575 144.600 109.855 ;
        RECT 0.055 97.755 144.320 98.575 ;
        RECT 0.055 85.775 144.600 97.755 ;
        RECT 0.055 84.955 144.320 85.775 ;
        RECT 0.055 73.675 144.600 84.955 ;
        RECT 0.055 72.855 144.320 73.675 ;
        RECT 0.055 60.875 144.600 72.855 ;
        RECT 0.055 60.055 144.320 60.875 ;
        RECT 0.055 48.775 144.600 60.055 ;
        RECT 0.055 47.955 144.320 48.775 ;
        RECT 0.055 35.975 144.600 47.955 ;
        RECT 0.055 35.155 144.320 35.975 ;
        RECT 0.055 23.875 144.600 35.155 ;
        RECT 0.055 23.055 144.320 23.875 ;
        RECT 0.055 12.850 144.600 23.055 ;
        RECT 0.055 12.030 144.320 12.850 ;
        RECT 0.055 11.850 144.600 12.030 ;
        RECT 0.055 11.030 144.320 11.850 ;
        RECT 0.055 10.850 144.600 11.030 ;
        RECT 0.055 10.030 144.320 10.850 ;
        RECT 0.055 9.850 144.600 10.030 ;
        RECT 0.055 9.030 144.320 9.850 ;
        RECT 0.055 8.850 144.600 9.030 ;
        RECT 0.055 8.030 144.320 8.850 ;
        RECT 0.055 7.850 144.600 8.030 ;
        RECT 0.055 7.030 144.320 7.850 ;
        RECT 0.055 6.850 144.600 7.030 ;
        RECT 0.055 6.030 144.320 6.850 ;
        RECT 0.055 5.850 144.600 6.030 ;
        RECT 0.055 5.030 144.320 5.850 ;
        RECT 0.055 4.850 144.600 5.030 ;
        RECT 0.055 4.030 144.320 4.850 ;
        RECT 0.055 3.850 144.600 4.030 ;
        RECT 0.055 3.030 144.320 3.850 ;
        RECT 0.055 2.850 144.600 3.030 ;
        RECT 0.055 2.030 144.320 2.850 ;
        RECT 0.055 1.850 144.600 2.030 ;
        RECT 0.055 1.030 144.320 1.850 ;
        RECT 0.055 0.130 144.600 1.030 ;
      LAYER met3 ;
        RECT 1.245 11.765 144.350 112.115 ;
        RECT 130.685 10.845 144.350 11.765 ;
        RECT 137.750 9.095 144.350 10.845 ;
        RECT 139.155 7.045 144.350 9.095 ;
        RECT 1.245 0.615 144.350 7.045 ;
  END
END rom_tvbgone_32k
END LIBRARY

